package yapp_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "/home/Raid_Al-Tamimi/Verification/Labs/Lab8/Task1_uvc/sv/yapp_packet.sv"
`include "/home/Raid_Al-Tamimi/Verification/Labs/Lab8/Task1_uvc/sv/yapp_tx_monitor.sv"
`include "/home/Raid_Al-Tamimi/Verification/Labs/Lab8/Task1_uvc/sv/yapp_tx_sequencer.sv"
`include "/home/Raid_Al-Tamimi/Verification/Labs/Lab8/Task1_uvc/sv/yapp_tx_seqs.sv"
`include "/home/Raid_Al-Tamimi/Verification/Labs/Lab8/Task1_uvc/sv/yapp_tx_driver.sv"
`include "/home/Raid_Al-Tamimi/Verification/Labs/Lab8/Task1_uvc/sv/yapp_tx_agent.sv"
`include "/home/Raid_Al-Tamimi/Verification/Labs/Lab8/Task1_uvc/tb/router_tb.sv"
`include "/home/Raid_Al-Tamimi/Verification/Labs/Lab8/Task1_uvc/tb/router_test_lib.sv"


endpackage